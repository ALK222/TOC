ENTITY nombre IS
    GENERIC (lista_de_parametros);
    PORT (
        A : IN BIT;
        B : OUT BIT);
END nombre;
