identificador : PROCESS (lista de sensibilidad)
BEGIN
    -- Sentencias secuenciales
    -- Sentencias condicionales
    -- Ecuaciones booleanas
END PROCESS; -- identificador
