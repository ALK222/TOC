id : FOR var IN rango LOOP
    list_of_statements
END LOOP id; -- id
