ENTITY F IS
    PORT (
        A, B : IN STD_LOGIC;
        Y : OUT STD_LOGIC);
END F;

ARCHITECTURE circuito OF F IS

    SIGNAL D, E : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL H : STD_LOGIC;

BEGIN

    -- Implementación del circuito

END circuito; -- circuito
