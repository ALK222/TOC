id : WHILE condition LOOP
    list_of_statements
END LOOP id; --id
