CASE expresion IS
    WHEN choice_1 => statements;
    WHEN choice_n => statemens;
    WHEN OTHERS => statemenst;
END CASE;
