PACKAGE nombre IS
    -- tipos personalizados
    -- constantes
    -- declaraciones de componentes
    -- funciones y procedimientos (SOLO declaraciones)
END nombre;

PACKAGE BODY nombre IS
    -- Funciones y procedimientos (cuerpo)
END nombre;
