id : LOOP
    list_of_statements
    -- Use exit statement to get ount
END LOOP id; -- id
