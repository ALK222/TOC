WITH id SELECT
    signal_name <= valor1 WHEN valor_id1,
    valor2 WHEN valor_id2,
    valori WHEN valor_idi,
    otro_valor WHEN OTHERS;
