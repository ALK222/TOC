ARCHITECTURE circuito OF nombre IS
    -- Signals
BEGIN
    -- Definición del circuito
END circuito; -- circuito
