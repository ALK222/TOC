signal_name <= valor_1 WHEN condition1 ELSE
    valor_2 WHEN condition2 ELSE
    valor_i WHEN condition1 ELSE
    otro_valor;
